`ifndef constants
`define constants


`typedef enum logic [6:0] {
    //Simple Fixed
    ADD_WORD = 7'd1;
    ADD_WORD_IMMEDIATE = 7'd2
    SUBTRACT_FROM_WORD = 7'd3
    SUBTRACT_FROM_IMMEDIATE= 7'd4
    ADD_EXTENDED = 7'd5
    CARRY_GENERATE = 7'd6
    SUBTRACT_FROM_EXTENDED = 7'd7
    BORROW_GENERATE = 7'd8
    ADD_HALFWORD= 7'd9
    ADD_HALFWORD_IMMEDIATE= 7'd10
    SUBTRACT_FROM_HALFWORD = 7'd11
    SUBTRACT_FROM_HALFWORD_IMMEDIATE = 7'd12
    COUNT_LEADING_ZEROS = 7'd13
    FORM_SELECT_MASK_FOR_HALFWORD = 7'd14
    FORM_SELECT_MARK_FOR_WORDS = 7'd15
    AND = 7'd16
    AND_WITH_COMPLEMENT = 7'd17
    AND_HALFWORD_IMMEDIATE = 7'd18
    AND_WORD_IMMEDIATE = 7'd19
    OR = 7'd20
    OR_WITH_COMPLEMENT = 7'd21
    OR_HALFWORD_IMMEDIATE= 7'd22
    OR_WORD_IMMEDIATE= 7'd23
    EXCLUSIVE_OR = 7'd24
    EXCLUSIVE_OR_HALFWORD_IMMEDIATE = 7'd25
    EXCLUSIVE_OR_WORD_IMMEDIATE = 7'd26
    NAND = 7'd27
    NOR = 7'd28
    COMPARE_EQUAL_HALFWORD = 7'd29
    COMPARE_EQUAL_HALFWORD_IMMEDIATE = 7'd30
    COMPARE_EQUAL_WORD = 7'd31
    COMPARE_EQUAL_WORD_IMMEDIATE = 7'd32
    COMPARE_GREATER_THAN_HALFWORD = 7'd33
    COMPARE_GREATER_THAN_HALFWORD_IMMEDIATE = 7'd34
    COMPARE_GREATER_THAN_WORD = 7'd35
    COMPARE_GREATER_THAN_WORD_IMMEDIATE = 7'd36
    COMPARE_LOGICAL_GREATER_THAN_HALFWORD = 7'd37
    COMPARE_LOGICAL_GREATER_THAN_HALFWORD_IMMEDIATE = 7'd38
    COMPARE_LOGICAL_GREATER_THAN_WORD = 7'd39
    COMPARE_LOGICAL_GREATER_THAN_WORD_IMMEDIATE = 7'd40
= 7'd41
= 7'd42
= 7'd43
= 7'd44
= 7'd45
= 7'd46
= 7'd47
= 7'd48
= 7'd49
= 7'd50
= 7'd51
= 7'd52
= 7'd53
= 7'd54
= 7'd55
= 7'd56
= 7'd57
= 7'd58
= 7'd59
= 7'd60
= 7'd61
= 7'd62
= 7'd63
= 7'd64
= 7'd65
= 7'd66
= 7'd67
= 7'd68
= 7'd69
= 7'd70
= 7'd71
= 7'd72
= 7'd73
= 7'd74
= 7'd75
= 7'd76
= 7'd77
= 7'd78
= 7'd79
= 7'd80
= 7'd81
= 7'd82
= 7'd83
= 7'd84
= 7'd85
= 7'd86
= 7'd87
= 7'd88
= 7'd89
= 7'd90

} internal_opcodes;

`endif 